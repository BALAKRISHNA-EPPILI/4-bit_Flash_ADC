* c:\ebalakrishna\fossee\esim\bala_priority_encoder\comp\comp.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/8/2022 12:52:09 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R2-Pad1_ vref vin Net-_X1-Pad4_ Net-_R2-Pad2_ Net-_R1-Pad1_ Net-_X1-Pad7_ ? lm_741		
v2  Net-_X1-Pad7_ GND 15		
v1  vin GND sine		
U2  vout plot_v1		
U1  vin plot_v1		
v4  GND Net-_X1-Pad4_ 15		
v3  vref GND 12		
U3  Net-_R1-Pad1_ vout adc_bridge_1		
R1  Net-_R1-Pad1_ GND 1k		
U4  vref plot_v1		
R2  Net-_R2-Pad1_ Net-_R2-Pad2_ 1k		

.end
